import zacore_common::*;

module zacore_decode_immediate #(

) (
    input inst_t inst,

    output w_t imm,
);

/* TODO */

endmodule
